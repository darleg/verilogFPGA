//NOT gate logic modeling
module NotGL(a,na);
input a;
output na;

not(na,a);
                
endmodule