module switchOn(output LED);

assign LED = 1;

endmodule