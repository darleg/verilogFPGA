module switchOff(output LED);

assign LED = 0;

endmodule